module register_8_bit(
	input logic CLK, Reset, Load, Shift_Enable, Shift_In,
	input logic [7:0] Data_In,
	output logic Shift_Out,
	output logic [7:0] Data_Out
);

	always_ff @ (posedge CLK)
	begin
	
	if(Reset)
		Data_Out <= 8'h0;
	else if(Load)
		Data_Out <= Data_In;
	else if(Shift_Enable)
		Data_Out <= {Shift_In, Data_Out[7:1]};
	end
	
	assign Shift_Out = Data_Out[0];
	
endmodule