module control_unit(
	input logic CLK, Reset, ClearA_LoadB, Execute, Register_B_Shift_Out,
	output logic Clear_Load, Shift, Load_XA, Subtract_Enable, Clear_Register
);

	enum logic [4:0] {start, load, add_0, shift_0,
											 add_1, shift_1,
											 add_2, shift_2,
											 add_3, shift_3,
											 add_4, shift_4,
											 add_5, shift_5,
											 add_6, shift_6,
											 add_7, shift_7,
							hold, check, restart} current_state, next_state;

	always_ff @ (posedge CLK or posedge Reset)
		begin
			if(Reset)
				current_state <= start;
			else
				current_state <= next_state;
		end
	
	always_comb
		begin
			next_state = current_state;
			
			unique case(current_state)
				
				start: 	if(ClearA_LoadB)
								next_state = load;
							
							else if(Execute)
								next_state = add_0;
				
				load: next_state = start;
				
				add_0:	next_state = shift_0;
				shift_0:	next_state = add_1;
				
				add_1:	next_state = shift_1;
				shift_1:	next_state = add_2;
				
				add_2:	next_state = shift_2;
				shift_2:	next_state = add_3;
				
				add_3:	next_state = shift_3;
				shift_3:	next_state = add_4;
				
				add_4:	next_state = shift_4;
				shift_4:	next_state = add_5;
				
				add_5:	next_state = shift_5;
				shift_5:	next_state = add_6;
				
				add_6:	next_state = shift_6;
				shift_6:	next_state = add_7;
				
				add_7:	next_state = shift_7;
				shift_7:	next_state = hold;
				
				hold:    if(~Execute)
								next_state = check;
				
				check:	if(Execute)
								next_state = restart;

				restart: next_state = add_0;
			endcase
		end

	always_comb
		begin
			case(current_state)
				
				start:
					begin
						Clear_Load = 1'b0;
						Shift = 1'b0;
						Load_XA = 1'b0;
						Subtract_Enable = 1'b0;
						Clear_Register = 1'b0;
					end
				
				load:
					begin
						Clear_Load = 1'b1;
						Shift = 1'b0;
						Load_XA = 1'b0;
						Subtract_Enable = 1'b0;
						Clear_Register = 1'b0;
					end
					
				add_0, add_1, add_2, add_3, add_4, add_5, add_6:
					begin
						Clear_Load = 1'b0;
						Shift = 1'b0;
						if(Register_B_Shift_Out)
							Load_XA = 1'b1;
						else
							Load_XA = 1'b0;
							Subtract_Enable = 1'b0;
							Clear_Register = 1'b0;
					end
				
				add_7:
					begin
						Clear_Load = 1'b0;
						Shift =1'b0;
						if(Register_B_Shift_Out)
							begin
								Load_XA = 1'b1;
								Subtract_Enable = 1'b1;
							end
						else
							begin
								Load_XA = 1'b0;
								Subtract_Enable <= 1'b0;
							end
						Clear_Register = 1'b0;
					end
				
				shift_0, shift_1, shift_2, shift_3, shift_4, shift_5, shift_6, shift_7:
					begin
						Clear_Load = 1'b0;
						Shift = 1'b1;
						Load_XA = 1'b0;
						Subtract_Enable = 1'b0;
						Clear_Register = 1'b0;
					end
				
				hold:
					begin
						Clear_Load <= 1'b0;
						Shift <= 1'b0;
						Load_XA <= 1'b0;
						Subtract_Enable = 1'b0;
						Clear_Register = 1'b0;
					end
					
				check:
					begin
						Clear_Load = 1'b0;
						Shift = 1'b0;
						Load_XA = 1'b0;
						Subtract_Enable = 1'b0;
						Clear_Register = 1'b0;
					end
				
				restart:
					begin
						Clear_Load = 1'b1;
						Shift = 1'b0;
						Load_XA = 1'b0;
						Subtract_Enable = 1'b0;
						Clear_Register = 1'b1;
					end
			endcase
		end

endmodule